`include "lib/defines.vh"
module ID(
    input wire clk,
    input wire rst,
    input wire [`StallBus-1:0] stall,
    
    output wire stallreq,

    input wire [`IF_TO_ID_WD-1:0] if_to_id_bus,//IF段传给ID段的数据，相当于IF_ID中间段模块

    input wire [31:0] inst_sram_rdata,//上一步中IF取到的指令

    input wire [`WB_TO_RF_WD-1:0] wb_to_rf_bus,//WB段传给ID段的数据

    output wire [`ID_TO_EX_WD-1:0] id_to_ex_bus,//ID段要传给EX段的数据，相当于ID_EX中间段

    output wire [`BR_WD-1:0] br_bus //跳转指令，传给IF段的
);

    reg [`IF_TO_ID_WD-1:0] if_to_id_bus_r;
    wire [31:0] inst;
    wire [31:0] id_pc;
    wire ce;
    //WB段回传数据
    wire wb_rf_we;
    wire [4:0] wb_rf_waddr;
    wire [31:0] wb_rf_wdata;

    always @ (posedge clk) begin//这一块实际上起到IF_ID模块的作用
        if (rst) begin
            if_to_id_bus_r <= `IF_TO_ID_WD'b0;        
        end else if (stall[1]==`Stop && stall[2]==`NoStop) begin
            if_to_id_bus_r <= `IF_TO_ID_WD'b0;//如果复位或者暂停的话就不要IF段传过来的数据了
        end else if (stall[1]==`NoStop) begin
            if_to_id_bus_r <= if_to_id_bus;
        end
    end
    
    assign inst = inst_sram_rdata;//inst就是上一步中IF取到的32位指令
    assign {//把IF_ID块解包
        ce,
        id_pc
    } = if_to_id_bus_r;
    assign {//把WB段回传数据解包
        wb_rf_we,
        wb_rf_waddr,
        wb_rf_wdata
    } = wb_to_rf_bus;
    
    //分解IF段取到的指令inst，划分为以下片段
    wire [5:0] opcode;
    wire [4:0] rs,rt,rd,sa;
    wire [5:0] func;
    wire [15:0] imm;
    wire [25:0] instr_index;
    wire [19:0] code;
    wire [4:0] base;
    wire [15:0] offset;
    wire [2:0] sel;
    assign opcode =       inst[31:26];
    assign rs =           inst[25:21];
    assign rt =           inst[20:16];
    assign rd =           inst[15:11];
    assign sa =           inst[10:6];
    assign func =         inst[5:0];
    assign imm =          inst[15:0];//立即数
    assign instr_index =  inst[25:0];
    assign code =         inst[25:6];
    assign base =         inst[25:21];
    assign offset =       inst[15:0];
    assign sel =          inst[2:0];

    wire [2:0] sel_alu_src1;
    wire [3:0] sel_alu_src2;
    wire [11:0] alu_op;

    wire data_ram_en;
    wire [3:0] data_ram_wen;
    
    wire rf_we;
    wire [4:0] rf_waddr;
    wire sel_rf_res;
    wire [2:0] sel_rf_dst;

    wire [31:0] rdata1, rdata2;

    regfile u_regfile(//对寄存器操作
    	.clk    (clk    ),
        .re1    (),//寄存器1是否可读
        .raddr1 (rs ),//读取的第一个寄存器rs
        .rdata1 (rdata1 ),//rs中读出来的数据
        .re2    (),//寄存器2是否可读
        .raddr2 (rt ),//读取的第二个寄存器rt
        .rdata2 (rdata2 ),//rt中读出来的数据
        .we     (wb_rf_we     ),//是否能写入寄存器
        .waddr  (wb_rf_waddr  ),//写入的寄存器地址
        .wdata  (wb_rf_wdata  )//写入的内容
    );

    wire inst_ori, inst_lui, inst_addiu, inst_beq;

    wire op_add, op_sub, op_slt, op_sltu;
    wire op_and, op_nor, op_or, op_xor;
    wire op_sll, op_srl, op_sra, op_lui;
    
    wire [63:0] op_d, func_d;
    decoder_6_64 u0_decoder_6_64(
    	.in  (opcode  ),
        .out (op_d )
    );

    decoder_6_64 u1_decoder_6_64(
    	.in  (func  ),
        .out (func_d )
    );
    
    wire [31:0] rs_d, rt_d, rd_d, sa_d;
    decoder_5_32 u0_decoder_5_32(
    	.in  (rs  ),
        .out (rs_d )
    );

    decoder_5_32 u1_decoder_5_32(
    	.in  (rt  ),
        .out (rt_d )
    );

    
    assign inst_ori     = op_d[6'b00_1101];//若opc是001101，则这个为1，代表译码得出是ori指令
    assign inst_lui     = op_d[6'b00_1111];//若opc是001111，则这个为1，代表译码得出是lui指令
    assign inst_addiu   = op_d[6'b00_1001];
    assign inst_beq     = op_d[6'b00_0100];



    // rs to reg1
    assign sel_alu_src1[0] = inst_ori | inst_addiu;

    // pc to reg1
    assign sel_alu_src1[1] = 1'b0;

    // sa_zero_extend to reg1
    assign sel_alu_src1[2] = 1'b0;

    
    // rt to reg2
    assign sel_alu_src2[0] = 1'b0;
    
    // imm_sign_extend to reg2
    assign sel_alu_src2[1] = inst_lui | inst_addiu;

    // 32'b8 to reg2
    assign sel_alu_src2[2] = 1'b0;

    // imm_zero_extend to reg2
    assign sel_alu_src2[3] = inst_ori;

    assign op_add = inst_addiu;
    assign op_sub = 1'b0;
    assign op_slt = 1'b0;
    assign op_sltu = 1'b0;
    assign op_and = 1'b0;
    assign op_nor = 1'b0;
    assign op_or = inst_ori;
    assign op_xor = 1'b0;
    assign op_sll = 1'b0;
    assign op_srl = 1'b0;
    assign op_sra = 1'b0;
    assign op_lui = inst_lui;

    //在下一步中，ALU算术逻辑单元要执行什么任务，对应的那一位就是1
    assign alu_op = {op_add, op_sub, op_slt, op_sltu,
                     op_and, op_nor, op_or, op_xor,
                     op_sll, op_srl, op_sra, op_lui};
    //这个alu_op会传给EX段


    // load and store enable
    assign data_ram_en = 1'b0;

    // write enable
    assign data_ram_wen = 1'b0;



    // regfile store enable
    assign rf_we = inst_ori | inst_lui | inst_addiu;



    // store in [rd]
    assign sel_rf_dst[0] = 1'b0;
    // store in [rt] 
    assign sel_rf_dst[1] = inst_ori | inst_lui | inst_addiu;
    // store in [31]
    assign sel_rf_dst[2] = 1'b0;

    // sel for regfile address
    assign rf_waddr = {5{sel_rf_dst[0]}} & rd 
                    | {5{sel_rf_dst[1]}} & rt
                    | {5{sel_rf_dst[2]}} & 32'd31;

    // 0 from alu_res ; 1 from ld_res
    assign sel_rf_res = 1'b0; 

    assign id_to_ex_bus = {
        id_pc,          // 158:127
        inst,           // 126:95
        alu_op,         // 94:83
        sel_alu_src1,   // 82:80
        sel_alu_src2,   // 79:76
        data_ram_en,    // 75
        data_ram_wen,   // 74:71
        rf_we,          // 70
        rf_waddr,       // 69:65
        sel_rf_res,     // 64
        rdata1,         // 63:32
        rdata2          // 31:0
    };

    //以下应该是beq相等转移指令的内容
    wire br_e;
    wire [31:0] br_addr;
    wire rs_eq_rt;//这个beq指令有用到
    wire rs_ge_z;//下面这四个都对应其它的跳转指令，让我们自己扩展的，比如这个应该是对应bgtz指令
    wire rs_gt_z;
    wire rs_le_z;
    wire rs_lt_z;
    wire [31:0] pc_plus_4;
    assign pc_plus_4 = id_pc + 32'h4;

    assign rs_eq_rt = (rdata1 == rdata2);//rs和rt的值是否相等？

    assign br_e = inst_beq & rs_eq_rt;//若确实是beq指令且rs和rt的值相等，那么可以跳转
    assign br_addr = inst_beq ? (pc_plus_4 + {{14{inst[15]}},inst[15:0],2'b0}) : 32'b0;
    //是beq指令，则跳转地址；否则跳转地址设为0
    assign br_bus = {
        br_e,
        br_addr
    };
    


endmodule